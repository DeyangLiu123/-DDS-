module rom(
	input clk,
    input[8:0] address, 
    output[11:0] data
);
	
	reg[11:0] r_data;
	
always @(posedge clk) begin
    case(address[7:0])
		8'd0:r_data<=12'b011111111111;
		8'd1:r_data<=12'b100000011000;
		8'd2:r_data<=12'b100000110001;
		8'd3:r_data<=12'b100001001010;
		8'd4:r_data<=12'b100001100011;
		8'd5:r_data<=12'b100001111100;
		8'd6:r_data<=12'b100010010101;
		8'd7:r_data<=12'b100010101110;
		8'd8:r_data<=12'b100011000111;
		8'd9:r_data<=12'b100011100000;
		8'd10:r_data<=12'b100011111001;
		8'd11:r_data<=12'b100100010010;
		8'd12:r_data<=12'b100100101011;
		8'd13:r_data<=12'b100101000100;
		8'd14:r_data<=12'b100101011100;
		8'd15:r_data<=12'b100101110101;
		8'd16:r_data<=12'b100110001110;
		8'd17:r_data<=12'b100110100110;
		8'd18:r_data<=12'b100110111111;
		8'd19:r_data<=12'b100111010111;
		8'd20:r_data<=12'b100111110000;
		8'd21:r_data<=12'b101000001000;
		8'd22:r_data<=12'b101000100000;
		8'd23:r_data<=12'b101000111001;
		8'd24:r_data<=12'b101001010001;
		8'd25:r_data<=12'b101001101001;
		8'd26:r_data<=12'b101010000001;
		8'd27:r_data<=12'b101010011000;
		8'd28:r_data<=12'b101010110000;
		8'd29:r_data<=12'b101011001000;
		8'd30:r_data<=12'b101011011111;
		8'd31:r_data<=12'b101011110111;
		8'd32:r_data<=12'b101100001110;
		8'd33:r_data<=12'b101100100101;
		8'd34:r_data<=12'b101100111100;
		8'd35:r_data<=12'b101101010011;
		8'd36:r_data<=12'b101101101010;
		8'd37:r_data<=12'b101110000000;
		8'd38:r_data<=12'b101110010111;
		8'd39:r_data<=12'b101110101101;
		8'd40:r_data<=12'b101111000011;
		8'd41:r_data<=12'b101111011010;
		8'd42:r_data<=12'b101111101111;
		8'd43:r_data<=12'b110000000101;
		8'd44:r_data<=12'b110000011011;
		8'd45:r_data<=12'b110000110000;
		8'd46:r_data<=12'b110001000110;
		8'd47:r_data<=12'b110001011011;
		8'd48:r_data<=12'b110001110000;
		8'd49:r_data<=12'b110010000101;
		8'd50:r_data<=12'b110010011001;
		8'd51:r_data<=12'b110010101110;
		8'd52:r_data<=12'b110011000010;
		8'd53:r_data<=12'b110011010110;
		8'd54:r_data<=12'b110011101010;
		8'd55:r_data<=12'b110011111110;
		8'd56:r_data<=12'b110100010001;
		8'd57:r_data<=12'b110100100100;
		8'd58:r_data<=12'b110100111000;
		8'd59:r_data<=12'b110101001010;
		8'd60:r_data<=12'b110101011101;
		8'd61:r_data<=12'b110101110000;
		8'd62:r_data<=12'b110110000010;
		8'd63:r_data<=12'b110110010100;
		8'd64:r_data<=12'b110110100110;
		8'd65:r_data<=12'b110110111000;
		8'd66:r_data<=12'b110111001001;
		8'd67:r_data<=12'b110111011010;
		8'd68:r_data<=12'b110111101011;
		8'd69:r_data<=12'b110111111100;
		8'd70:r_data<=12'b111000001101;
		8'd71:r_data<=12'b111000011101;
		8'd72:r_data<=12'b111000101101;
		8'd73:r_data<=12'b111000111101;
		8'd74:r_data<=12'b111001001100;
		8'd75:r_data<=12'b111001011100;
		8'd76:r_data<=12'b111001101011;
		8'd77:r_data<=12'b111001111010;
		8'd78:r_data<=12'b111010001000;
		8'd79:r_data<=12'b111010010110;
		8'd80:r_data<=12'b111010100101;
		8'd81:r_data<=12'b111010110010;
		8'd82:r_data<=12'b111011000000;
		8'd83:r_data<=12'b111011001101;
		8'd84:r_data<=12'b111011011010;
		8'd85:r_data<=12'b111011100111;
		8'd86:r_data<=12'b111011110100;
		8'd87:r_data<=12'b111100000000;
		8'd88:r_data<=12'b111100001100;
		8'd89:r_data<=12'b111100010111;
		8'd90:r_data<=12'b111100100011;
		8'd91:r_data<=12'b111100101110;
		8'd92:r_data<=12'b111100111001;
		8'd93:r_data<=12'b111101000100;
		8'd94:r_data<=12'b111101001110;
		8'd95:r_data<=12'b111101011000;
		8'd96:r_data<=12'b111101100010;
		8'd97:r_data<=12'b111101101011;
		8'd98:r_data<=12'b111101110100;
		8'd99:r_data<=12'b111101111101;
		8'd100:r_data<=12'b111110000110;
		8'd101:r_data<=12'b111110001110;
		8'd102:r_data<=12'b111110010110;
		8'd103:r_data<=12'b111110011110;
		8'd104:r_data<=12'b111110100101;
		8'd105:r_data<=12'b111110101101;
		8'd106:r_data<=12'b111110110011;
		8'd107:r_data<=12'b111110111010;
		8'd108:r_data<=12'b111111000000;
		8'd109:r_data<=12'b111111000110;
		8'd110:r_data<=12'b111111001100;
		8'd111:r_data<=12'b111111010001;
		8'd112:r_data<=12'b111111010110;
		8'd113:r_data<=12'b111111011011;
		8'd114:r_data<=12'b111111011111;
		8'd115:r_data<=12'b111111100100;
		8'd116:r_data<=12'b111111100111;
		8'd117:r_data<=12'b111111101011;
		8'd118:r_data<=12'b111111101110;
		8'd119:r_data<=12'b111111110001;
		8'd120:r_data<=12'b111111110100;
		8'd121:r_data<=12'b111111110110;
		8'd122:r_data<=12'b111111111000;
		8'd123:r_data<=12'b111111111010;
		8'd124:r_data<=12'b111111111011;
		8'd125:r_data<=12'b111111111100;
		8'd126:r_data<=12'b111111111101;
		8'd127:r_data<=12'b111111111101;
		8'd128:r_data<=12'b111111111110;
		8'd129:r_data<=12'b111111111101;
		8'd130:r_data<=12'b111111111101;
		8'd131:r_data<=12'b111111111100;
		8'd132:r_data<=12'b111111111011;
		8'd133:r_data<=12'b111111111010;
		8'd134:r_data<=12'b111111111000;
		8'd135:r_data<=12'b111111110110;
		8'd136:r_data<=12'b111111110100;
		8'd137:r_data<=12'b111111110001;
		8'd138:r_data<=12'b111111101110;
		8'd139:r_data<=12'b111111101011;
		8'd140:r_data<=12'b111111100111;
		8'd141:r_data<=12'b111111100100;
		8'd142:r_data<=12'b111111011111;
		8'd143:r_data<=12'b111111011011;
		8'd144:r_data<=12'b111111010110;
		8'd145:r_data<=12'b111111010001;
		8'd146:r_data<=12'b111111001100;
		8'd147:r_data<=12'b111111000110;
		8'd148:r_data<=12'b111111000000;
		8'd149:r_data<=12'b111110111010;
		8'd150:r_data<=12'b111110110011;
		8'd151:r_data<=12'b111110101101;
		8'd152:r_data<=12'b111110100101;
		8'd153:r_data<=12'b111110011110;
		8'd154:r_data<=12'b111110010110;
		8'd155:r_data<=12'b111110001110;
		8'd156:r_data<=12'b111110000110;
		8'd157:r_data<=12'b111101111101;
		8'd158:r_data<=12'b111101110100;
		8'd159:r_data<=12'b111101101011;
		8'd160:r_data<=12'b111101100010;
		8'd161:r_data<=12'b111101011000;
		8'd162:r_data<=12'b111101001110;
		8'd163:r_data<=12'b111101000100;
		8'd164:r_data<=12'b111100111001;
		8'd165:r_data<=12'b111100101110;
		8'd166:r_data<=12'b111100100011;
		8'd167:r_data<=12'b111100010111;
		8'd168:r_data<=12'b111100001100;
		8'd169:r_data<=12'b111100000000;
		8'd170:r_data<=12'b111011110100;
		8'd171:r_data<=12'b111011100111;
		8'd172:r_data<=12'b111011011010;
		8'd173:r_data<=12'b111011001101;
		8'd174:r_data<=12'b111011000000;
		8'd175:r_data<=12'b111010110010;
		8'd176:r_data<=12'b111010100101;
		8'd177:r_data<=12'b111010010110;
		8'd178:r_data<=12'b111010001000;
		8'd179:r_data<=12'b111001111010;
		8'd180:r_data<=12'b111001101011;
		8'd181:r_data<=12'b111001011100;
		8'd182:r_data<=12'b111001001100;
		8'd183:r_data<=12'b111000111101;
		8'd184:r_data<=12'b111000101101;
		8'd185:r_data<=12'b111000011101;
		8'd186:r_data<=12'b111000001101;
		8'd187:r_data<=12'b110111111100;
		8'd188:r_data<=12'b110111101011;
		8'd189:r_data<=12'b110111011010;
		8'd190:r_data<=12'b110111001001;
		8'd191:r_data<=12'b110110111000;
		8'd192:r_data<=12'b110110100110;
		8'd193:r_data<=12'b110110010100;
		8'd194:r_data<=12'b110110000010;
		8'd195:r_data<=12'b110101110000;
		8'd196:r_data<=12'b110101011101;
		8'd197:r_data<=12'b110101001010;
		8'd198:r_data<=12'b110100111000;
		8'd199:r_data<=12'b110100100100;
		8'd200:r_data<=12'b110100010001;
		8'd201:r_data<=12'b110011111110;
		8'd202:r_data<=12'b110011101010;
		8'd203:r_data<=12'b110011010110;
		8'd204:r_data<=12'b110011000010;
		8'd205:r_data<=12'b110010101110;
		8'd206:r_data<=12'b110010011001;
		8'd207:r_data<=12'b110010000101;
		8'd208:r_data<=12'b110001110000;
		8'd209:r_data<=12'b110001011011;
		8'd210:r_data<=12'b110001000110;
		8'd211:r_data<=12'b110000110000;
		8'd212:r_data<=12'b110000011011;
		8'd213:r_data<=12'b110000000101;
		8'd214:r_data<=12'b101111101111;
		8'd215:r_data<=12'b101111011010;
		8'd216:r_data<=12'b101111000011;
		8'd217:r_data<=12'b101110101101;
		8'd218:r_data<=12'b101110010111;
		8'd219:r_data<=12'b101110000000;
		8'd220:r_data<=12'b101101101010;
		8'd221:r_data<=12'b101101010011;
		8'd222:r_data<=12'b101100111100;
		8'd223:r_data<=12'b101100100101;
		8'd224:r_data<=12'b101100001110;
		8'd225:r_data<=12'b101011110111;
		8'd226:r_data<=12'b101011011111;
		8'd227:r_data<=12'b101011001000;
		8'd228:r_data<=12'b101010110000;
		8'd229:r_data<=12'b101010011000;
		8'd230:r_data<=12'b101010000001;
		8'd231:r_data<=12'b101001101001;
		8'd232:r_data<=12'b101001010001;
		8'd233:r_data<=12'b101000111001;
		8'd234:r_data<=12'b101000100000;
		8'd235:r_data<=12'b101000001000;
		8'd236:r_data<=12'b100111110000;
		8'd237:r_data<=12'b100111010111;
		8'd238:r_data<=12'b100110111111;
		8'd239:r_data<=12'b100110100110;
		8'd240:r_data<=12'b100110001110;
		8'd241:r_data<=12'b100101110101;
		8'd242:r_data<=12'b100101011100;
		8'd243:r_data<=12'b100101000100;
		8'd244:r_data<=12'b100100101011;
		8'd245:r_data<=12'b100100010010;
		8'd246:r_data<=12'b100011111001;
		8'd247:r_data<=12'b100011100000;
		8'd248:r_data<=12'b100011000111;
		8'd249:r_data<=12'b100010101110;
		8'd250:r_data<=12'b100010010101;
		8'd251:r_data<=12'b100001111100;
		8'd252:r_data<=12'b100001100011;
		8'd253:r_data<=12'b100001001010;
		8'd254:r_data<=12'b100000110001;
		8'd255:r_data<=12'b100000011000;

    endcase
end

	assign data = address[8] ? 12'b111111111110 - r_data : r_data; 

endmodule